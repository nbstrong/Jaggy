library ieee;
use ieee.std_logic_1164.all;

-- Arithmetic Logic Unit
entity arith_log_unit is
	port (datain1, datain2: in std_logic_vector(31 downto 0);
		dataout: out std_logic_vector(31 downto 0));
end arith_log_unit;

architecture struct of arith_log_unit is
begin
end struct;